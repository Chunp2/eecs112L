module  processorTb;
//----------------------Processor-----------------------
reg ref_clk;
reg reset;

Processor L1(
	.ref_clk(ref_clk),
	.reset(reset)
	);

initial
	 begin 
	reset=1; 

	#10 
	reset=0;
	ref_clk = 0; 
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10 
	reset=0;
	ref_clk = 0; 
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10 
	reset=0;
	ref_clk = 0; 
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10 
	reset=0;
	ref_clk = 0; 
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10 
	reset=0;
	ref_clk = 0; 
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
	#10;
	ref_clk = 0; 
	reset=0;
	#10; 
	ref_clk = 1; 
	reset=0;
end 
endmodule
